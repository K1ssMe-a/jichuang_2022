`define DATA_WIDTH 8
`define DATA_ZERO  8'b0
`define COEFF_ZERO 10'b0
`define MUTI_ZERO  17'b0

`define LCDI_IDLE   3'd0
`define LCDI_STATE1 3'd1
`define LCDI_STATE2 3'd2
`define LCDI_STATE3 3'd3
`define LCDI_STATE4 3'd4
`define LCDI_STATE5 3'd5
`define LCDI_STATE6 3'd6        
